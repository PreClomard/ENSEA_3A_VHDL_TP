-------------------------------------------------------------------------------------------
-- Testbench pour DCPT_M avec deux compteurs
-------------------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tst_dcpt_m is
end tst_dcpt_m;

architecture tst_dcpt_m_arch of tst_dcpt_m is
  constant CLK_PERIOD : time := 10 ns;
  constant M : integer := 2;  -- Exemple : M=4 pour le premier compteur

  -- Signaux pour le premier compteur (M bits)
  signal ENABLE_M : STD_LOGIC := '0';
  signal UD_M     : STD_LOGIC := '0';
  signal RESET_M  : STD_LOGIC := '0';
  signal CPTR_M   : STD_LOGIC_VECTOR(M-1 downto 0);

  -- Signaux pour le deuxieme compteur (8 bits)
  signal ENABLE_8 : STD_LOGIC := '0';
  signal UD_8     : STD_LOGIC := '0';
  signal RESET_8  : STD_LOGIC := '0';
  signal CPTR_8   : STD_LOGIC_VECTOR(7 downto 0);

  -- Signal d'horloge commun
  signal CLK : STD_LOGIC := '0';

  -- Composant DCPT_M
  component DCPT_M
    generic (
      M : integer
    );
    port (
      ENABLE : in  STD_LOGIC;
      UD     : in  STD_LOGIC;
      RESET  : in  STD_LOGIC;
      CLK    : in  STD_LOGIC;
      CPTR   : out STD_LOGIC_VECTOR(M-1 downto 0)
    );
  end component;

begin
  -- Instance du premier compteur (M bits)
  uut_M: DCPT_M
    generic map (M => M)
    port map (
      ENABLE => ENABLE_M,
      UD     => UD_M,
      RESET  => RESET_M,
      CLK    => CLK,
      CPTR   => CPTR_M
    );

  -- Instance du deuxieme compteur (8 bits)
  uut_8: DCPT_M
    generic map (M => 8)
    port map (
      ENABLE => ENABLE_8,
      UD     => UD_8,
      RESET  => RESET_8,
      CLK    => CLK,
      CPTR   => CPTR_8
    );

  -- Generation d'horloge commune
  CLK_process: process
  begin
    CLK <= '0';
    wait for CLK_PERIOD/2;
    CLK <= '1';
    wait for CLK_PERIOD/2;
  end process;

  -- Stimulus pour le premier compteur (M bits)
  stimulus_M: process
  begin
    -- R�initialisation
    RESET_M <= '1';
    wait for 20 ns;
    RESET_M <= '0';

    -- Activation du comptage
    ENABLE_M <= '1';
    UD_M <= '1';  -- Mode compteur
    wait for 200 ns;

    -- Changer en mode deecompteur
    UD_M <= '0';
    wait for 200 ns;

    -- Desactiver le comptage/decomptage
    ENABLE_M <= '0';
    wait;
  end process;

  -- Stimulus pour le deuxieme compteur (8 bits)
  stimulus_8: process
  begin
    -- Reinitialisation
    RESET_8 <= '1';
    wait for 20 ns;
    RESET_8 <= '0';

    -- Activation du comptage
    ENABLE_8 <= '1';
    UD_8 <= '1';  -- Mode compteur
    wait for 200 ns;

    -- Changer en mode decompteur
    UD_8 <= '0';
    wait for 200 ns;

    -- Desactiver le comptage/deecomptage
    ENABLE_8 <= '0';
    wait;
  end process;

end tst_dcpt_m_arch;
