library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity complement_a_2_tb is
end complement_a_2_tb;

architecture Behavioral of complement_a_2_tb is
    constant N : integer := 8; -- 8 bits par mot

    signal nombre  : STD_LOGIC_VECTOR(N-1 downto 0);
    signal sortie  : STD_LOGIC_VECTOR(N-1 downto 0);

begin
    -- Instanciation
    uut: entity work.complement_a_2
        generic map (N => N)
        port map (
            nombre   => nombre,
            sortie  => sortie
        );

    -- Stimuli
    stim_proc: process
    begin

        nombre <= "10101010"; wait for 20 ns;
	nombre <= "11111111"; wait for 20 ns;
	nombre <= "11110000"; wait for 20 ns;
        -- Fin de simulation
        wait;
    end process;
end Behavioral;

