library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.FIFO_Component.all;

entity FastSlow is
  generic (
    M : integer := 4  -- Par d�faut, M=4 pour une FIFO de 16 mots
  );
  port (
    CLK      : in  STD_LOGIC;
    Incwrite : in  STD_LOGIC;
    Incread  : in  STD_LOGIC;
    Reset_in    : in STD_LOGIC;
    Fast     : out STD_LOGIC;  -- '1' si le nombre de mots dans la FIFO est < 2^(M-2)
    Slow     : out STD_LOGIC   -- '1' si le nombre de mots dans la FIFO est >= 2^M - 2^(M-2)
  );
end FastSlow;

architecture Behavioral of FastSlow is
  signal counter_value : STD_LOGIC_VECTOR(M-1 downto 0) := (others => '0');

begin
    write_counter_inst: DCPT_M
    generic map (M => M)
    port map (
      ENABLE  => '1',
      UD      => Incwrite,
      RESET   => Reset_in,
      CLK     => CLK,
      CPTR    => counter_value
    );

  -- Logique pour g�n�rer les signaux Fast et Slow
  Fast <= '1' when to_integer(unsigned(counter_value)) < 2**(M-2) else '0';
  Slow <= '1' when to_integer(unsigned(counter_value)) >= (2**M - 2**(M-2)) else '0';

end Behavioral;

