library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package FIFO_Component is

-- Declaration du composant DCPT_M (Compteur/Decompteur M bits)
  component DCPT_M
    generic (
      M : integer := 8
    );
    port (
      ENABLE : in  STD_LOGIC; 
      UD     : in  STD_LOGIC; 
      RESET  : in  STD_LOGIC; 
      CLK    : in  STD_LOGIC; 
      CPTR   : out STD_LOGIC_VECTOR(M-1 downto 0) 
    );
  end component;

  -- Declaration du composant GENHL (Generateur d'horloge de lecture)
  component GENHL
    generic (
      Div : integer := 200  -- Valeur de division
    );
    port (
      RESET   : in  STD_LOGIC;
      CLK     : in  STD_LOGIC;
      ENREAD  : out STD_LOGIC;
      ENWRITE : out STD_LOGIC
    );
  end component;

  -- Declaration du composant RAM
  component RAM
    generic (
      M : integer := 4;  
      N : integer := 8  
    );
    port (
      CS_n  : in  STD_LOGIC; 
      RW_n  : in  STD_LOGIC; 
      OE    : in  STD_LOGIC;  
      Adr   : in  STD_LOGIC_VECTOR(M-1 downto 0);
      Din   : in  STD_LOGIC_VECTOR(N-1 downto 0);
      Dout  : out STD_LOGIC_VECTOR(N-1 downto 0)
    );
  end component;

  -- Declaration du composant MUX_M2to1 (Multiplexeur M x 2 vers 1)
component MUX_M2to1
  generic (
    M : integer := 4  -- Taille des bus d'entr�e
  );
  port (
    A   : in  STD_LOGIC_VECTOR(M-1 downto 0);
    B   : in  STD_LOGIC_VECTOR(M-1 downto 0);
    SEL : in  STD_LOGIC;
    Y   : out STD_LOGIC_VECTOR(M-1 downto 0)
  );
end component;

  -- Declaration du composant GENADR (Generateur d'adresse)
  component GENADR
    generic (
      M : integer := 4 
    );
    port (
      RESET    : in  STD_LOGIC;
      CLK      : in  STD_LOGIC;
      incread  : in  STD_LOGIC;
      incwrite : in  STD_LOGIC;
      selread  : in  STD_LOGIC;
      Adrg     : out STD_LOGIC_VECTOR(M-1 downto 0)
    );
  end component;

  -- Declaration du composant FASTSLOW
  component FASTSLOW
    generic (
      M : integer := 4
    );
    port (
      RESET    : in  STD_LOGIC;
      CLK      : in  STD_LOGIC;
      incread  : in  STD_LOGIC;
      incwrite : in  STD_LOGIC;
      fast     : out STD_LOGIC;
      slow     : out STD_LOGIC
    );
  end component;

  -- Declaration du composant complement_a_2
  component complement_a_2
    generic (
      N : natural := 8
    );
    port (
      nombre : in  std_logic_vector(N-1 downto 0);
      sortie : out std_logic_vector(N-1 downto 0)
    );
  end component;

  -- Declaration du composant Reg_N (Registre N bits)
  component Reg_N
    generic (
      N : integer := 8
    );
    port (
      RESET : in  STD_LOGIC;
      CLK   : in  STD_LOGIC;
      D     : in  STD_LOGIC_VECTOR(N-1 downto 0);
      Q     : out STD_LOGIC_VECTOR(N-1 downto 0)
    );
  end component;

  -- Declaration du composant SEQUENCEUR
  component sequenceur
    port (
      enwrite, enread, clk, reset, req : in  STD_LOGIC; 
      acq, rw_n, oe, incwrite, incread, hl, selread, cs_n : out STD_LOGIC
    );
  end component;

end package FIFO_Component;
